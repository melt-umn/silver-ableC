grammar edu:umn:cs:melt:exts:silver:ableC:concretesyntax;

exports edu:umn:cs:melt:exts:silver:ableC:concretesyntax:quotation;
exports edu:umn:cs:melt:exts:silver:ableC:concretesyntax:antiquotation;

exports edu:umn:cs:melt:ableC:concretesyntax;
exports edu:umn:cs:melt:ableC:concretesyntax:construction;
